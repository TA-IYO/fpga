module fnd_top(

);


endmodule